--
--	Package File Template
--
--	Purpose: This package defines supplemental types, subtypes, 
--		 constants, and functions 
--
--   To use any of the example code shown below, uncomment the lines and modify as necessary
--

library IEEE;
use IEEE.STD_LOGIC_1164.all;

package MIPS_package is

-- type <new_type> is
--  record
--    <type_name>        : std_logic_vector( 7 downto 0);
--    <type_name>        : std_logic;
-- end record;
--
-- Declare constants
--
-- constant <constant_name>		: time := <time_unit> ns;
-- constant <constant_name>		: integer := <value;
--
-- Declare functions and procedure
--
-- function <function_name>  (signal <signal_name> : in <type_declaration>) return <type_declaration>;
-- procedure <procedure_name> (<type_declaration> <constant_name>	: in <type_declaration>);
--
subtype bus32 is std_logic_vector(31 downto 0);
subtype bus16 is std_logic_vector(15 downto 0);
subtype bus7 is std_logic_vector	(6 downto 0);
subtype bus6 is std_logic_vector (5 downto 0);
subtype bus5 is std_logic_vector (4 downto 0);
subtype bus4 is std_logic_vector (3 downto 0);
subtype bus2 is std_logic_vector (1 downto 0);
subtype bus1 is std_logic;

COMPONENT instruction_memory
  PORT (
    clka : IN STD_LOGIC;
    addra : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
  );
END COMPONENT;

COMPONENT register_bank
PORT(
	read_address1 : IN std_logic_vector(4 downto 0);
	read_address2 : IN std_logic_vector(4 downto 0);
	write_address : IN std_logic_vector(4 downto 0);
	data_in : IN std_logic_vector(31 downto 0);
	write_en : IN std_logic;
	clock : IN std_logic;          
	data_out1 : OUT std_logic_vector(31 downto 0);
	data_out2 : OUT std_logic_vector(31 downto 0)
	);
END COMPONENT;

COMPONENT ALU
	PORT(
		ALU_op : IN std_logic_vector(3 downto 0);
		input1 : IN std_logic_vector(31 downto 0);
		input2 : IN std_logic_vector(31 downto 0);          
		output : OUT std_logic_vector(31 downto 0);
		zero : OUT std_logic
		);
END COMPONENT;

COMPONENT data_mem
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
  );
END COMPONENT;

type micro_code is 
	record
	branch: bus1;  -- '1' If it's branch instruction
	jump:   bus1;  -- '1' If it's jump instruction
	reg_op1: bus1; -- '1' If register1 needs to be readed
	reg_op2: bus1; -- '1' If register2 needs to be readed
	imm_sign: bus1;  -- '1' If immediate operand is sign extended
	reg_dest_select: bus2; -- what type of destiny register, rt"00" or rd"01", or ra"11"
	reg_write: bus1; -- '1' If the operation involves a register write
	R_or_I: bus1;   -- whether ALU operates on two registers '0' or register and immediate '1'
	mem_op: bus1;  -- '1' If the operation involves memory access
	mem_write: bus1;  -- '1' If the memory operation is a write
	ALU_op: bus4;  -- ALU control signal
	reg_result_select: bus2;  -- what to be written in to register. "00" ALU output, "01" data memory output, "11" PC+4
end record;	

type micro_code_table is array (0 to 127) of micro_code;
-- ** stands for instructions that exist in MIPS but not implemented in our design
-- NOP: not an operation
constant my_mips_code: micro_code_table :=
(
--b,  j, r1, r2, sig, des, rw, I, mo, mw, ALU_op,A/M/P
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --0   
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --1    
('0','1','0','0','0',"00",'0','0','0','0',"1111","00"),  --2   j   
('0','1','0','0','0',"11",'1','0','0','0',"1111","11"),	--3   jal  
('1','0','1','1','1',"00",'0','0','0','0',"0110","00"),  --4   beq 
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --5   bne  **
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --6   blez **
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --7   bgtz **
('0','0','1','0','1',"00",'1','1','0','0',"0010","00"),  --8   addi :no exception raised
('0','0','1','0','0',"00",'1','1','0','0',"0010","00"),  --9   addiu :no exception, no sign extension (different from actual MIPS)
('0','0','1','0','1',"00",'1','1','0','0',"0111","00"),  --10  slti  
('0','0','1','0','0',"00",'1','1','0','0',"0111","00"),	--11  sltiu  
('0','0','1','0','1',"00",'1','1','0','0',"0000","00"),  --12  andi
('0','0','1','0','1',"00",'1','1','0','0',"0001","00"),  --13  ori
('0','0','1','0','1',"00",'1','1','0','0',"0100","00"),  --14  xori
('0','0','0','0','0',"00",'1','1','0','0',"1111","00"),  --15	lui
--b,  j, r1, r2, sig, des, rw, I, mo, mw, ALU_op,A/M/P
('0','0','0','0','0',"10",'0','0','0','0',"1111","00"),  --16  Speicial test register
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --17
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --18
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),	--19
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --20
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --21
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --22
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --23
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --24
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --25
('0','1','0','0','0',"00",'0','0','0','0',"1111","00"),  --26 
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),	--27 
('1','0','1','1','1',"00",'0','0','0','0',"1111","00"),  --28
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --29
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --30 
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --31  
--b,  j, r1, r2, sig, des, rw, I, mo, mw, ALU_op,A/M/P
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --32  lb **
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --33	lh **
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --34	lwl **
('0','0','1','0','1',"00",'1','1','1','0',"0010","01"),	--35  lw
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --36  lbu **
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --37  lhu **
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --38 	lwr **
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --39  NOP
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --40  sb **
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --41	sh **
('0','1','0','0','0',"00",'0','0','0','0',"1111","00"),  --42 	swl **
('0','0','1','1','1',"00",'0','1','1','1',"0010","00"),	--43	sw
--b,  j, r1, r2, sig, des, rw, I, mo, mw, ALU_op,A/M/P
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --44
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --45
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --46	swr **
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --47	cache **
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --48	ll**
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --49	lwc1**
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --50 	lwc2**
('0','0','0','0','0',"00",'0','0','0','0',"1111","11"),	--51  pref**
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --52
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --53	ldc1**
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --54 	ldc2**
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --55
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --56	sc**
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --57	swc1**
--b,  j, r1, r2, sig, des, rw, I, mo, mw, ALU_op,A/M/P
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --58 	swc2**
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),	--59 
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --60
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --61	sdc1**
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --62 	sdc2**
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),	--63
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --64  sll(in this implementation this instr will be fetched when all '0')
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --65
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --66 
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),	--67 
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --68
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --69
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --70 
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),	--71
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --72
--b,  j, r1, r2, sig, des, rw, I, mo, mw, ALU_op,A/M/P
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --73
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --74 
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),	--75 
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --76
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --77
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --78 
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),	--79
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --80
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --81
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --82
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),	--83 
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --84
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --85
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --86 
--b,  j, r1, r2, sig, des, rw, I, mo, mw, ALU_op,A/M/P
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),	--87
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --88
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --89
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --90 
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),	--91 
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --92
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --93
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --94 
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),	--95
('0','0','1','1','0',"01",'1','0','0','0',"0010","00"),  --96	add
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --97	addu** (no point implementing this when no exception supported)
('0','0','1','1','0',"01",'1','0','0','0',"0110","00"),  --98 	sub
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),	--99 	subu** same reason as above
('0','0','1','1','0',"01",'1','0','0','0',"0000","00"),  --100 and
('0','0','1','1','0',"01",'1','0','0','0',"0001","00"),  --101 or
('0','0','1','1','0',"01",'1','0','0','0',"0100","00"),  --102 xor
--b,  j, r1, r2, sig, des, rw, I, mo, mw, ALU_op,A/M/P
('0','0','1','1','0',"01",'1','0','0','0',"0011","00"),	--103 nor
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --104
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --105
('0','0','1','1','0',"01",'1','0','0','0',"0111","00"),  --106 slt
('0','0','0','0','0',"11",'0','0','0','0',"1111","11"),	--107 sltu** same reason as above
('1','0','1','1','1',"00",'0','0','0','0',"1111","00"),  --108
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --109
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --110 
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),	--111
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --112
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --113
('0','1','0','0','0',"00",'0','0','0','0',"1111","00"),  --114
('0','0','0','0','0',"11",'0','0','0','0',"1111","11"),	--115 
--b,  j, r1, r2, sig, des, rw, I, mo, mw, ALU_op,A/M/P
('1','0','1','1','1',"00",'0','0','0','0',"1111","00"),  --116
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --117
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --118 
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),	--119
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --120
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --121
('0','1','0','0','0',"00",'0','0','0','0',"1111","00"),  --122 
('0','0','0','0','0',"11",'0','0','0','0',"1111","11"),	--123 
('1','0','1','1','1',"00",'0','0','0','0',"1111","00"),  --124
('0','0','0','0','0',"00",'0','0','0','0',"1101","00"),  --125
('0','0','0','0','0',"00",'0','0','0','0',"1111","00"),  --126
('0','0','0','0','0',"00",'0','0','0','0',"1111","00")	--127
);

type bank_type is array (1 to 31) of bus32;
	
end MIPS_package;

package body MIPS_package is

---- Example 1
--  function <function_name>  (signal <signal_name> : in <type_declaration>  ) return <type_declaration> is
--    variable <variable_name>     : <type_declaration>;
--  begin
--    <variable_name> := <signal_name> xor <signal_name>;
--    return <variable_name>; 
--  end <function_name>;

---- Example 2
--  function <function_name>  (signal <signal_name> : in <type_declaration>;
--                         signal <signal_name>   : in <type_declaration>  ) return <type_declaration> is
--  begin
--    if (<signal_name> = '1') then
--      return <signal_name>;
--    else
--      return 'Z';
--    end if;
--  end <function_name>;

---- Procedure Example
--  procedure <procedure_name>  (<type_declaration> <constant_name>  : in <type_declaration>) is
--    
--  begin
--    
--  end <procedure_name>;
 
end MIPS_package;
